module DUT(
);
endmodule;
