module DUT(
    input write_port,
    input [127:0] write_quad_port,
    input write_array_port [0:127],
    input [127:0] write_quad_array_port [0:127],
    input reg write_reg_port,
    input wire write_wire_port
);

endmodule;
